--------------------------------------------
-- Author:            Miquel Saula
-- Last modification: 3/08/2020
--------------------------------------------

Library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

entity execution_module is
    generic (
        -- System
        SA: integer:= 32;
        SD: integer:= 32;
        SX: integer:= 17;
        SB: integer:= 5;

        -- Instruction
        IO: integer:= 4;
        IX: integer:= 2;
        IY: integer:= 11;

        -- Floating Point
        FD: integer:= 32;
        FM: integer:= 23;
        FE: integer:= 8;

        BC: integer:= 8
    );
    port (
        clk: in std_logic;
        reset: in std_logic;
        EXE_Stall: in std_logic;

        -- Connexions amb el IDM
        A: in std_logic_vector(SD-1 downto 0);
        B: in std_logic_vector(SD-1 downto 0);
        Af: in std_logic_vector(SD-1 downto 0);
        Bf: in std_logic_vector(SD-1 downto 0);

        InstructionToExecute: in std_logic_vector(SX-1 downto 0);
        RD: in std_logic_vector(SB-1 downto 0);

        BPIDQ: out std_logic_vector(SD-1 downto 0);
        BPIDIFP: out std_logic;
        BPIDNFI: out std_logic;

        BPEXERD: out std_logic_vector(SB-1 downto 0);
        BPEXEIFP: out std_logic;
        BPEXENFI: out std_logic;

        -- Conexions amb el MEM
        InstructionExecuted: out std_logic_vector(SX-1 downto 0);
        ALUOut: out std_logic_vector(SD-1 downto 0);
        SMDR: out std_logic_vector(SD-1 downto 0);
        cond: out std_logic;

        -- Altres connexions
        ALUNotReady: out std_logic;
        ret: out std_logic;
        LIFOout: in std_logic_vector(SD-1 downto 0);

        -- OoOE Bus
        ACK0: in std_logic;
        Q0: out std_logic_vector(FD-1 downto 0);
        RD0: out std_logic_vector(SB-1 downto 0);
        END0: out std_logic;
        IFP0: out std_logic;

        ACK1: in std_logic;
        Q1: out std_logic_vector(FD-1 downto 0);
        RD1: out std_logic_vector(SB-1 downto 0);
        END1: out std_logic;
        IFP1: out std_logic;

        ACK2: in std_logic;
        Q2: out std_logic_vector(FD-1 downto 0);
        RD2: out std_logic_vector(SB-1 downto 0);
        END2: out std_logic;
        IFP2: out std_logic;

        ACK3: in std_logic;
        Q3: out std_logic_vector(FD-1 downto 0);
        RD3: out std_logic_vector(SB-1 downto 0);
        END3: out std_logic;
        IFP3: out std_logic;

        ACK4: in std_logic;
        Q4: out std_logic_vector(FD-1 downto 0);
        RD4: out std_logic_vector(SB-1 downto 0);
        END4: out std_logic;
        IFP4: out std_logic;

        ACK5: in std_logic;
        Q5: out std_logic_vector(FD-1 downto 0);
        RD5: out std_logic_vector(SB-1 downto 0);
        END5: out std_logic;
        IFP5: out std_logic;

        ACK6: in std_logic;
        Q6: out std_logic_vector(FD-1 downto 0);
        RD6: out std_logic_vector(SB-1 downto 0);
        END6: out std_logic;
        IFP6: out std_logic;

        ACK7: in std_logic;
        Q7: out std_logic_vector(FD-1 downto 0);
        RD7: out std_logic_vector(SB-1 downto 0);
        END7: out std_logic;
        IFP7: out std_logic
	);
end execution_module;

architecture a of execution_module is

    component fpu is
        generic (
            -- System
            SX: integer:= 17;
            SB: integer:= 5;

            -- Instruction
            IO: integer:= 4;
            IX: integer:= 2;
            IY: integer:= 11;

            -- Floating Point
            FD: integer:= 32;
            FM: integer:= 23;
            FE: integer:= 8;

            BC: integer:= 8
        );
        port (
            clk: in std_logic;
            reset: in std_logic;
            EXE_Stall: in std_logic;

            InstructionToExecute: in std_logic_vector(SX-1 downto 0);

            A: in std_logic_vector(SD-1 downto 0);
            B: in std_logic_vector(SD-1 downto 0);

            C: out std_logic_vector(SD-1 downto 0);

            FPUNotReady: out std_logic;

            RDin: in std_logic_vector(SB-1 downto 0);
            IsFP: in std_logic;

            -- OoOE Bus
            ACK0: in std_logic;
            Q0: out std_logic_vector(FD-1 downto 0);
            RD0: out std_logic_vector(SB-1 downto 0);
            END0: out std_logic;
            IFP0: out std_logic;

            ACK1: in std_logic;
            Q1: out std_logic_vector(FD-1 downto 0);
            RD1: out std_logic_vector(SB-1 downto 0);
            END1: out std_logic;
            IFP1: out std_logic;

            ACK2: in std_logic;
            Q2: out std_logic_vector(FD-1 downto 0);
            RD2: out std_logic_vector(SB-1 downto 0);
            END2: out std_logic;
            IFP2: out std_logic;

            ACK3: in std_logic;
            Q3: out std_logic_vector(FD-1 downto 0);
            RD3: out std_logic_vector(SB-1 downto 0);
            END3: out std_logic;
            IFP3: out std_logic;

            ACK4: in std_logic;
            Q4: out std_logic_vector(FD-1 downto 0);
            RD4: out std_logic_vector(SB-1 downto 0);
            END4: out std_logic;
            IFP4: out std_logic;

            ACK5: in std_logic;
            Q5: out std_logic_vector(FD-1 downto 0);
            RD5: out std_logic_vector(SB-1 downto 0);
            END5: out std_logic;
            IFP5: out std_logic;

            ACK6: in std_logic;
            Q6: out std_logic_vector(FD-1 downto 0);
            RD6: out std_logic_vector(SB-1 downto 0);
            END6: out std_logic;
            IFP6: out std_logic;

            ACK7: in std_logic;
            Q7: out std_logic_vector(FD-1 downto 0);
            RD7: out std_logic_vector(SB-1 downto 0);
            END7: out std_logic;
            IFP7: out std_logic
    	);
    end component;

    component int2sevseg is
        port (
            input: in std_logic_vector(SD-1 downto 0);
            output: out std_logic_vector(SD-1 downto 0)
        );
    end component;

    constant all_ones: std_logic_vector(SD-1 downto 0) := (others => '1');
    constant all_zero: std_logic_vector(SD-1 downto 0) := (others => '0');

    signal C: std_logic_vector(SD-1 downto 0) := (others => '0');

    signal Ai: integer := 0;
    signal Bi: integer := 0;
    signal Ci: integer := 0;

    signal opcode: std_logic_vector(IO-1 downto 0) := (others => '0');
    signal flags: std_logic_vector(IX-1 downto 0) := (others => '0');
    signal flags2: std_logic_vector(IY-1 downto 0) := (others => '0');

    signal shiftAux: std_logic_vector(SD-1 downto 0) := (others => '0');
    signal sevsegAux: std_logic_vector(SD-1 downto 0) := (others => '0');
    signal FPUOut: std_logic_vector(FD-1 downto 0) := (others => '0');

    signal isfp: std_logic;

    signal InstructionExecutedAux: std_logic_vector(SX-1 downto 0);

begin

    FPUU: fpu
    generic map (
        SX => SX,
        SB => SB,

        IO => IO,
        IX => IX,
        IY => IY,

        FD => FD,
        FM => FM,
        FE => FE,

        BC => BC
    ) port map (
        clk => clk,
        reset => reset,
        EXE_Stall => EXE_Stall,
        InstructionToExecute => InstructionToExecute,
        A => A,
        B => B,
        C => FPUOut,
        FPUNotReady => ALUNotReady,
        RDin => RD,
        IsFP => isfp,
        ACK0 => ACK0,
        Q0 => Q0,
        RD0 => RD0,
        END0 => END0,
        IFP0 => IFP0,
        ACK1 => ACK1,
        Q1 => Q1,
        RD1 => RD1,
        END1 => END1,
        IFP1 => IFP1,
        ACK2 => ACK2,
        Q2 => Q2,
        RD2 => RD2,
        END2 => END2,
        IFP2 => IFP2,
        ACK3 => ACK3,
        Q3 => Q3,
        RD3 => RD3,
        END3 => END3,
        IFP3 => IFP3,
        ACK4 => ACK4,
        Q4 => Q4,
        RD4 => RD4,
        END4 => END4,
        IFP4 => IFP4,
        ACK5 => ACK5,
        Q5 => Q5,
        RD5 => RD5,
        END5 => END5,
        IFP5 => IFP5,
        ACK6 => ACK6,
        Q6 => Q6,
        RD6 => RD6,
        END6 => END6,
        IFP6 => IFP6,
        ACK7 => ACK7,
        Q7 => Q7,
        RD7 => RD7,
        END7 => END7,
        IFP7 => IFP7
    );

    I2SS: int2sevseg
    port map (
        input => A,
        output => sevsegAux
    );

    isfp <= '1' when (opcode = "0000" and flags = "10") or (opcode = "0100" and flags = "01") else '0';

    opcode <= InstructionToExecute(IO-1 downto 0);
    flags <= InstructionToExecute((IO+IX)-1 downto IO);
    flags2 <= InstructionToExecute((IO+IX+IY)-1 downto (IO+IX));

    Ai <= to_integer(unsigned(A));
    Bi <= to_integer(unsigned(B));

    Ci <=
        Ai + Bi when opcode = "0000" and flags = "00" and flags2 = "00000000000" else
        Ai + Bi when opcode = "0000" and flags = "01" else
        Ai - Bi when opcode = "0000" and flags = "00" and flags2 = "00000000001" else
        Ai * Bi when opcode = "0000" and flags = "00" and flags2 = "00000000010" else
        Ai / Bi when opcode = "0000" and flags = "00" and flags2 = "00000000011" else
        to_integer(unsigned(A AND B)) when opcode = "0001" and flags = "00" and flags2 = "00000000000" else
        to_integer(unsigned(A OR B))  when opcode = "0001" and flags = "00" and flags2 = "00000000001" else
        to_integer(unsigned(A XOR B)) when opcode = "0001" and flags = "00" and flags2 = "00000000010" else
        to_integer(unsigned(NOT A)) +1 when opcode = "0001" and flags = "00" and flags2 = "00000000011" else
        to_integer(unsigned(NOT A))    when opcode = "0001" and flags = "00" and flags2 = "00000000100" else
        to_integer(unsigned(sevsegAux)) when opcode = "1111" else
        to_integer(unsigned(B(15 downto 0) & A(15 downto 0))) when opcode = "0010" and flags = "00" else
        to_integer(unsigned(A(31 downto 16) & B(15 downto 0))) when opcode = "0010" and flags = "01" else
        to_integer(unsigned(shiftAux)) when opcode = "0011" else
        to_integer(unsigned(all_ones)) when Ai = Bi and opcode = "0101" and flags = "00" and flags2 = "00000000000" else
        to_integer(unsigned(all_zero)) when (not (Ai = Bi)) and opcode = "0101" and flags = "00" and flags2 = "00000000000" else
        to_integer(unsigned(all_ones)) when Ai > Bi and opcode = "0101" and flags = "00" and flags2 = "00000000001" else
        to_integer(unsigned(all_zero)) when (not (Ai > Bi)) and opcode = "0101" and flags = "00" and flags2 = "00000000001" else
        to_integer(unsigned(all_ones)) when Ai < Bi and opcode = "0101" and flags = "00" and flags2 = "00000000010" else
        to_integer(unsigned(all_zero)) when (not (Ai < Bi)) and opcode = "0101" and flags = "00" and flags2 = "00000000010" else
        Ai + Bi when opcode = "1101" else
        Ai + Bi when opcode = "1100" and flags = "00" else
        Ai + Bi when opcode = "1100" and flags = "01" else
        to_integer(unsigned(LIFOout)) +4 when opcode = "1100" and flags = "10" else
        Ai + Bi when opcode = "0111" or opcode = "1000" or opcode = "0110" else
        to_integer(unsigned(FPUOut)) when (((opcode = "0000") and (flags = "10")) or ((opcode = "0101") and (flags = "10"))) or (opcode = "0100") else
        to_integer(unsigned(all_zero));

    C <= std_logic_vector(to_signed(Ci, SD));

    BPIDQ <= C;
    BPIDIFP <= '1' when ((opcode = "0100") and (flags = "01")) or
                ((opcode = "0000") and (flags = "10")) else '0';-- or
                --((opcode = "0101") and (flags = "10") and (flags2 = "00000000001")) or
                --((opcode = "1101") and (flags = "10")) else '0';
    BPEXEIFP <= '1' when ((InstructionExecutedAux(IO-1 downto 0) = "0100") and (InstructionExecutedAux(IO+IX-1 downto IO) = "00")) or
                ((InstructionExecutedAux(IO-1 downto 0) = "0000") and (InstructionExecutedAux(IO+IX-1 downto IO) = "10")) else '0';-- or
                --((InstructionExecutedAux(IO-1 downto 0) = "0101") and (InstructionExecutedAux(IO+IX-1 downto IO) = "10") and (InstructionExecutedAux(IO+IX+IY-1 downto IO+IX) = "00000000001")) or
                --((InstructionExecutedAux(IO-1 downto 0) = "1101") and (InstructionExecutedAux(IO+IX-1 downto IO) = "10")) else '0';

    BPIDNFI <= '1' when (opcode = "0000") and (flags = "10") and (flags2 = "00000000011") else '0';
    BPEXENFI <= '1' when (InstructionExecutedAux(IO-1 downto 0) = "0000") and (InstructionExecutedAux(IO+IX-1 downto IO) = "10") and (InstructionExecutedAux(IO+IX+IY-1 downto IO+IX) = "00000000011") else '0';

    ret <= '1' when InstructionToExecute(IO-1 downto 0) = "1100" and InstructionToExecute((IO+IX)-1 downto IO) = "10" else '0';

    InstructionExecuted <= InstructionExecutedAux;

    updateOutputs: process(clk)
    begin
        if (clk = '1' and EXE_Stall = '0') then
            if (opcode = "1100" and flags = "01") then SMDR <= B;
            else SMDR <= Bf; end if;

            InstructionExecutedAux <= InstructionToExecute;
            ALUOut <= C;

            BPEXERD <= RD;

            if (Af = Bf) then cond <= '1';
            else cond <= '0'; end if;
        end if;
    end process;

    performShiftOperation: process(Ai, Bi, opcode, flags, flags2)
    begin
        if (opcode = "0011") then
            if (Bi >= 32) then
                shiftAux <= (others => '0'); -- 0
            elsif (Bi < 0) then
                shiftAux <= (others => '1'); -- error
            else
                if (flags = "00") then
                    shiftAux(SD-1 downto Bi) <= A((SD-1) - Bi downto 0);
                    shiftAux(Bi-1 downto 0) <= (others => '0');
                elsif (flags = "01") then
                    shiftAux(SD - Bi -1 downto 0) <= A((SD-1) downto Bi);
                    if (flags2 = "00000000000") then
                        shiftAux((SD-1) downto SD - Bi) <= (others => '0');
                    elsif (flags2 = "00000000001") then
                        shiftAux((SD-1) downto SD - Bi) <= (others => A((SD-1)));
                    end if;
                end if;
            end if;
        end if;
    end process;

end a;
